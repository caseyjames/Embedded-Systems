// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// Revision Information:
// 05Feb10              Production Release Version 3.0
// SVN Revision Information:
// SVN $Revision: 12344 $
// SVN $Date: 2010-02-27 21:59:30 -0800 (Sat, 27 Feb 2010) $
`timescale 1ns/1ps
module
CAPB3O
(
input
[
15
:
0
]
CAPB3I,
input
[
31
:
0
]
PRDATAS0,
input
[
31
:
0
]
PRDATAS1,
input
[
31
:
0
]
PRDATAS2,
input
[
31
:
0
]
PRDATAS3,
input
[
31
:
0
]
PRDATAS4,
input
[
31
:
0
]
PRDATAS5,
input
[
31
:
0
]
PRDATAS6,
input
[
31
:
0
]
PRDATAS7,
input
[
31
:
0
]
PRDATAS8,
input
[
31
:
0
]
PRDATAS9,
input
[
31
:
0
]
PRDATAS10,
input
[
31
:
0
]
PRDATAS11,
input
[
31
:
0
]
PRDATAS12,
input
[
31
:
0
]
PRDATAS13,
input
[
31
:
0
]
PRDATAS14,
input
[
31
:
0
]
PRDATAS15,
input
[
15
:
0
]
CAPB3l,
input
[
15
:
0
]
CAPB3OI,
output
wire
PREADY,
output
wire
PSLVERR,
output
wire
[
31
:
0
]
PRDATA
)
;
localparam
[
3
:
0
]
CAPB3II
=
4
'b
0000
;
localparam
[
3
:
0
]
CAPB3lI
=
4
'b
0001
;
localparam
[
3
:
0
]
CAPB3Ol
=
4
'b
0010
;
localparam
[
3
:
0
]
CAPB3Il
=
4
'b
0011
;
localparam
[
3
:
0
]
CAPB3ll
=
4
'b
0100
;
localparam
[
3
:
0
]
CAPB3O0
=
4
'b
0101
;
localparam
[
3
:
0
]
CAPB3I0
=
4
'b
0110
;
localparam
[
3
:
0
]
CAPB3l0
=
4
'b
0111
;
localparam
[
3
:
0
]
CAPB3O1
=
4
'b
1000
;
localparam
[
3
:
0
]
CAPB3I1
=
4
'b
1001
;
localparam
[
3
:
0
]
CAPB3l1
=
4
'b
1010
;
localparam
[
3
:
0
]
CAPB3OOI
=
4
'b
1011
;
localparam
[
3
:
0
]
CAPB3IOI
=
4
'b
1100
;
localparam
[
3
:
0
]
CAPB3lOI
=
4
'b
1101
;
localparam
[
3
:
0
]
CAPB3OII
=
4
'b
1110
;
localparam
[
3
:
0
]
CAPB3III
=
4
'b
1111
;
reg
CAPB3lII
;
reg
CAPB3OlI
;
reg
[
31
:
0
]
CAPB3IlI
;
wire
[
3
:
0
]
CAPB3llI
;
wire
[
31
:
0
]
CAPB3O0I
;
assign
CAPB3O0I
=
32
'b
0
;
assign
CAPB3llI
[
3
]
=
CAPB3I
[
15
]
|
CAPB3I
[
14
]
|
CAPB3I
[
13
]
|
CAPB3I
[
12
]
|
CAPB3I
[
11
]
|
CAPB3I
[
10
]
|
CAPB3I
[
9
]
|
CAPB3I
[
8
]
;
assign
CAPB3llI
[
2
]
=
CAPB3I
[
15
]
|
CAPB3I
[
14
]
|
CAPB3I
[
13
]
|
CAPB3I
[
12
]
|
CAPB3I
[
7
]
|
CAPB3I
[
6
]
|
CAPB3I
[
5
]
|
CAPB3I
[
4
]
;
assign
CAPB3llI
[
1
]
=
CAPB3I
[
15
]
|
CAPB3I
[
14
]
|
CAPB3I
[
11
]
|
CAPB3I
[
10
]
|
CAPB3I
[
7
]
|
CAPB3I
[
6
]
|
CAPB3I
[
3
]
|
CAPB3I
[
2
]
;
assign
CAPB3llI
[
0
]
=
CAPB3I
[
15
]
|
CAPB3I
[
13
]
|
CAPB3I
[
11
]
|
CAPB3I
[
9
]
|
CAPB3I
[
7
]
|
CAPB3I
[
5
]
|
CAPB3I
[
3
]
|
CAPB3I
[
1
]
;
always
@(*)
begin
case
(
CAPB3llI
)
CAPB3II
:
if
(
CAPB3I
[
0
]
)
CAPB3IlI
[
31
:
0
]
=
PRDATAS0
[
31
:
0
]
;
else
CAPB3IlI
[
31
:
0
]
=
CAPB3O0I
[
31
:
0
]
;
CAPB3lI
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS1
[
31
:
0
]
;
CAPB3Ol
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS2
[
31
:
0
]
;
CAPB3Il
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS3
[
31
:
0
]
;
CAPB3ll
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS4
[
31
:
0
]
;
CAPB3O0
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS5
[
31
:
0
]
;
CAPB3I0
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS6
[
31
:
0
]
;
CAPB3l0
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS7
[
31
:
0
]
;
CAPB3O1
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS8
[
31
:
0
]
;
CAPB3I1
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS9
[
31
:
0
]
;
CAPB3l1
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS10
[
31
:
0
]
;
CAPB3OOI
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS11
[
31
:
0
]
;
CAPB3IOI
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS12
[
31
:
0
]
;
CAPB3lOI
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS13
[
31
:
0
]
;
CAPB3OII
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS14
[
31
:
0
]
;
CAPB3III
:
CAPB3IlI
[
31
:
0
]
=
PRDATAS15
[
31
:
0
]
;
default
:
CAPB3IlI
[
31
:
0
]
=
CAPB3O0I
[
31
:
0
]
;
endcase
end
always
@(*)
begin
case
(
CAPB3llI
)
CAPB3II
:
if
(
CAPB3I
[
0
]
)
CAPB3lII
=
CAPB3l
[
0
]
;
else
CAPB3lII
=
1
'b
1
;
CAPB3lI
:
CAPB3lII
=
CAPB3l
[
1
]
;
CAPB3Ol
:
CAPB3lII
=
CAPB3l
[
2
]
;
CAPB3Il
:
CAPB3lII
=
CAPB3l
[
3
]
;
CAPB3ll
:
CAPB3lII
=
CAPB3l
[
4
]
;
CAPB3O0
:
CAPB3lII
=
CAPB3l
[
5
]
;
CAPB3I0
:
CAPB3lII
=
CAPB3l
[
6
]
;
CAPB3l0
:
CAPB3lII
=
CAPB3l
[
7
]
;
CAPB3O1
:
CAPB3lII
=
CAPB3l
[
8
]
;
CAPB3I1
:
CAPB3lII
=
CAPB3l
[
9
]
;
CAPB3l1
:
CAPB3lII
=
CAPB3l
[
10
]
;
CAPB3OOI
:
CAPB3lII
=
CAPB3l
[
11
]
;
CAPB3IOI
:
CAPB3lII
=
CAPB3l
[
12
]
;
CAPB3lOI
:
CAPB3lII
=
CAPB3l
[
13
]
;
CAPB3OII
:
CAPB3lII
=
CAPB3l
[
14
]
;
CAPB3III
:
CAPB3lII
=
CAPB3l
[
15
]
;
default
:
CAPB3lII
=
1
'b
1
;
endcase
end
always
@(*)
begin
case
(
CAPB3llI
)
CAPB3II
:
if
(
CAPB3I
[
0
]
)
CAPB3OlI
=
CAPB3OI
[
0
]
;
else
CAPB3OlI
=
1
'b
0
;
CAPB3lI
:
CAPB3OlI
=
CAPB3OI
[
1
]
;
CAPB3Ol
:
CAPB3OlI
=
CAPB3OI
[
2
]
;
CAPB3Il
:
CAPB3OlI
=
CAPB3OI
[
3
]
;
CAPB3ll
:
CAPB3OlI
=
CAPB3OI
[
4
]
;
CAPB3O0
:
CAPB3OlI
=
CAPB3OI
[
5
]
;
CAPB3I0
:
CAPB3OlI
=
CAPB3OI
[
6
]
;
CAPB3l0
:
CAPB3OlI
=
CAPB3OI
[
7
]
;
CAPB3O1
:
CAPB3OlI
=
CAPB3OI
[
8
]
;
CAPB3I1
:
CAPB3OlI
=
CAPB3OI
[
9
]
;
CAPB3l1
:
CAPB3OlI
=
CAPB3OI
[
10
]
;
CAPB3OOI
:
CAPB3OlI
=
CAPB3OI
[
11
]
;
CAPB3IOI
:
CAPB3OlI
=
CAPB3OI
[
12
]
;
CAPB3lOI
:
CAPB3OlI
=
CAPB3OI
[
13
]
;
CAPB3OII
:
CAPB3OlI
=
CAPB3OI
[
14
]
;
CAPB3III
:
CAPB3OlI
=
CAPB3OI
[
15
]
;
default
:
CAPB3OlI
=
1
'b
0
;
endcase
end
assign
PREADY
=
CAPB3lII
;
assign
PSLVERR
=
CAPB3OlI
;
assign
PRDATA
=
CAPB3IlI
[
31
:
0
]
;
endmodule
